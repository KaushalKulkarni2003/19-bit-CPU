module PC_Adder(
    input [18:0] a,
    input [18:0] b,
    output [18:0] c
);

assign c= a + b;

endmodule